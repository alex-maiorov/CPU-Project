
typedef enum logic [3:0] {CONTROL_S, MEMORY_S, PC_S, ALU_S} systembus_mux_t;


module control(
input logic [31:0] 



endmodule
