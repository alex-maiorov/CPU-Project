module mul(a,
b,
clk,
signctl,
dout
)

endmodule

